library verilog;
use verilog.vl_types.all;
entity CPU_TB is
    generic(
        R0              : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        R1              : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        R2              : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        R3              : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        OP_LDW          : vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        OP_STW          : vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        OP_ADDI         : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        OP_BR           : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        OP_BLT          : vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        OP_BEQ          : vl_logic_vector(5 downto 0) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        OP_R            : vl_logic_vector(5 downto 0) := (Hi1, Hi1, Hi1, Hi0, Hi1, Hi0);
        OP_CALL         : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        OPX_ADD         : vl_logic_vector(10 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        OPX_SUB         : vl_logic_vector(10 downto 0) := (Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDR            : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BR_ADDR         : vl_logic_vector(15 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        LOAD_R1         : vl_logic_vector(31 downto 0);
        LOAD_R2         : vl_logic_vector(31 downto 0);
        STORE_R1        : vl_logic_vector(31 downto 0);
        ADDI_R1         : vl_logic_vector(31 downto 0);
        ADD_R1R2        : vl_logic_vector(31 downto 0);
        SUB_R1R2        : vl_logic_vector(31 downto 0);
        BR_START        : vl_logic_vector(31 downto 0);
        BR_R0R1         : vl_logic_vector(31 downto 0);
        CALL0           : vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of R0 : constant is 2;
    attribute mti_svvh_generic_type of R1 : constant is 2;
    attribute mti_svvh_generic_type of R2 : constant is 2;
    attribute mti_svvh_generic_type of R3 : constant is 2;
    attribute mti_svvh_generic_type of OP_LDW : constant is 2;
    attribute mti_svvh_generic_type of OP_STW : constant is 2;
    attribute mti_svvh_generic_type of OP_ADDI : constant is 2;
    attribute mti_svvh_generic_type of OP_BR : constant is 2;
    attribute mti_svvh_generic_type of OP_BLT : constant is 2;
    attribute mti_svvh_generic_type of OP_BEQ : constant is 2;
    attribute mti_svvh_generic_type of OP_R : constant is 2;
    attribute mti_svvh_generic_type of OP_CALL : constant is 2;
    attribute mti_svvh_generic_type of OPX_ADD : constant is 2;
    attribute mti_svvh_generic_type of OPX_SUB : constant is 2;
    attribute mti_svvh_generic_type of ADDR : constant is 2;
    attribute mti_svvh_generic_type of BR_ADDR : constant is 2;
    attribute mti_svvh_generic_type of LOAD_R1 : constant is 4;
    attribute mti_svvh_generic_type of LOAD_R2 : constant is 4;
    attribute mti_svvh_generic_type of STORE_R1 : constant is 4;
    attribute mti_svvh_generic_type of ADDI_R1 : constant is 4;
    attribute mti_svvh_generic_type of ADD_R1R2 : constant is 4;
    attribute mti_svvh_generic_type of SUB_R1R2 : constant is 4;
    attribute mti_svvh_generic_type of BR_START : constant is 4;
    attribute mti_svvh_generic_type of BR_R0R1 : constant is 4;
    attribute mti_svvh_generic_type of CALL0 : constant is 4;
end CPU_TB;
