module control(
    iClk, nRst, iPC,
    PC_en, IR_en, MDR_en, MAR_en,
    RF_Write,
    ALU_op,
    MAR_Select, ALUB_Select, AddrC_Select, PCA_Select,
    PC_Select, C_Select
);



endmodule
