module ha(
    a,
    b,
    sum,
    cout
);


input reg 
