module DE2_VGA (
    
);
    
endmodule