library verilog;
use verilog.vl_types.all;
entity ADDER_TB is
end ADDER_TB;
