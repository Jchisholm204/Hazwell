package charString is

    type characterString is array ( 0 to 31 ) of std_logic_vector(7 downto 0);

end package charString;

package body charString IS
end package body charString;