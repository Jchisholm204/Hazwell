library verilog;
use verilog.vl_types.all;
entity mux_using_assign_TB is
end mux_using_assign_TB;
