library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity top is
    port();
end entity;

architecture rtl of top is

begin

end architecture;