c1_inst : c1 PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);
