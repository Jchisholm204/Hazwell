entity test is
end entity;

architecture sim of test is
begin

	process is
		begin
		wait;
		end process;
end architecture;
